/**
 * PET Clone - Open hardware implementation of the Commodore PET
 * by Daniel Lehenbauer and contributors.
 * 
 * https://github.com/DLehenbauer/commodore-pet-clone
 *
 * To the extent possible under law, I, Daniel Lehenbauer, have waived all
 * copyright and related or neighboring rights to this project. This work is
 * published from the United States.
 *
 * @copyright CC0 http://creativecommons.org/publicdomain/zero/1.0/
 * @author Daniel Lehenbauer <DLehenbauer@users.noreply.github.com> and contributors
 */

// Implements core of SPI Mode 0 transfers in a controller/peripheral agnostic way.
 module spi #(
    parameter DATA_WIDTH = 8
) (
    // SPI bus signals (see https://www.oshwa.org/a-resolution-to-redefine-spi-signal-names/)
    input  logic spi_cs_ni,             // (CS)  Chip Select (active low)
    input  logic spi_sck_i,             // (SCK) Serial Clock
    input  logic spi_sd_i,              // (SDI) Serial Data In (rx)
    output logic spi_sd_o,              // (SDO) Serial Data Out (tx)
    
    // Relevant WB bus signals in SCK domain.
    input  logic [DATA_WIDTH-1:0] data_i,     // Data to transmit.  Captured on falling edge of CS_N and
                                              // falling edge of SCK for LSB.

    output logic [DATA_WIDTH-1:0] data_o,     // Data received.  Shifted in from SDO on each positive edge of SCK.
    
    output logic                  strobe_o    // Asserted on rising SCK when 'data_o' is valid.  The next 'data_i'
                                              // is captured on the following negative SCK edege.
);
    logic [$clog2(DATA_WIDTH-1)-1:0] bits_remaining = DATA_WIDTH-1;

    initial begin
        strobe_o <= '0;
    end

    logic [DATA_WIDTH-1:0] rx_buffer_d, rx_buffer_q;
    assign rx_buffer_d = { rx_buffer_q[DATA_WIDTH-2:0], spi_sd_i };

    logic [DATA_WIDTH-1:0] tx_buffer_q;
    logic preload = 1'b1;

    logic spi_sd_q;
    assign spi_sd_o = preload
        ? data_i[DATA_WIDTH-1]
        : spi_sd_q;
    
    wire msb = bits_remaining == DATA_WIDTH-1;
    wire lsb = bits_remaining == '0;

    always_ff @(posedge spi_cs_ni or posedge spi_sck_i) begin
        if (spi_cs_ni) begin
            // Deasserting 'spi_cs_ni' indicates the transfer has ended.
            bits_remaining <= DATA_WIDTH-1;
            rx_buffer_q    <= 'x;
            tx_buffer_q    <= 'x;
            strobe_o       <= '0;
        end else begin
            // SDI is valid on positive edge of SCK.
            rx_buffer_q <= rx_buffer_d;

            if (msb) tx_buffer_q    <= data_i;
            if (lsb) data_o         <= rx_buffer_d;

            strobe_o         <= lsb;
            bits_remaining <= bits_remaining - 1'b1;
        end
    end

    always_ff @(posedge spi_cs_ni or negedge spi_sck_i) begin
        if (spi_cs_ni) begin
            preload     <= 1'b1;
        end else begin
            spi_sd_q    <= tx_buffer_q[bits_remaining];
            preload     <= msb;
        end
    end
endmodule
